// Buffer in Verilog

module buffer(
	input A,
	output Y
);

assign Y = A;

endmodule
